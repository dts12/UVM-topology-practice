interface my_interface (input logic clock);

endinterface:my_interface